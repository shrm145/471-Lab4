library verilog;
use verilog.vl_types.all;
entity zeroFlag_testbench is
end zeroFlag_testbench;
