library verilog;
use verilog.vl_types.all;
entity controls_testbench is
end controls_testbench;
