library verilog;
use verilog.vl_types.all;
entity mux2_1_5Bit_testbench is
end mux2_1_5Bit_testbench;
