library verilog;
use verilog.vl_types.all;
entity decoder5x32_testbench is
end decoder5x32_testbench;
