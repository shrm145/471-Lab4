library verilog;
use verilog.vl_types.all;
entity nor32Bit_testbench is
end nor32Bit_testbench;
