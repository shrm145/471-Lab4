library verilog;
use verilog.vl_types.all;
entity calcSltu_testbench is
end calcSltu_testbench;
