library verilog;
use verilog.vl_types.all;
entity mux16_1_testbench is
end mux16_1_testbench;
